module main;
  initial $print_rust("hii");
endmodule