module main;
  initial $test1(42);
endmodule