module main;
  initial $bitvec(10'b1010101111);
endmodule